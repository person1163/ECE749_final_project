//----------------------------------------------------------------------
// Created with uvmf_gen version 2023.4_2
//----------------------------------------------------------------------
// pragma uvmf custom header begin
// pragma uvmf custom header end
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//
// DESCRIPTION: This package contains test level parameters
//
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//


package lc3_parameters_pkg;

  import uvmf_base_pkg_hdl::*;

  // pragma uvmf custom package_imports_additional begin 
  // pragma uvmf custom package_imports_additional end


  // These parameters are used to uniquely identify each interface.  The monitor_bfm and
  // driver_bfm are placed into and retrieved from the uvm_config_db using these string 
  // names as the field_name. The parameter is also used to enable transaction viewing 
  // from the command line for selected interfaces using the UVM command line processing.
  parameter string fetch_fetch_in_agent_BFM  = "fetch_fetch_in_agent_BFM"; /* [0] */
  parameter string fetch_fetch_out_agent_BFM  = "fetch_fetch_out_agent_BFM"; /* [1] */
  parameter string memaccess_memaccess_in_agent_BFM  = "memaccess_memaccess_in_agent_BFM"; /* [2] */
  parameter string memaccess_memaccess_out_agent_BFM  = "memaccess_memaccess_out_agent_BFM"; /* [3] */
  parameter string control_control_in_agent_BFM  = "control_control_in_agent_BFM"; /* [4] */
  parameter string control_control_out_agent_BFM  = "control_control_out_agent_BFM"; /* [5] */
  parameter string imem_agent_BFM  = "imem_agent_BFM"; /* [6] */
  parameter string dmem_agent_BFM  = "dmem_agent_BFM"; /* [7] */

  // pragma uvmf custom package_item_additional begin
  // pragma uvmf custom package_item_additional end

endpackage

// pragma uvmf custom external begin
// pragma uvmf custom external end


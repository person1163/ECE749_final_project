package decode_test_pkg;
    import uvm_pkg::*;
    import decode_in_pkg::*;
    import decode_out_pkg::*;
    import decode_env_pkg::*;
    import lc3_prediction_pkg::*;
    `include "uvm_macros.svh"
    `include "src/test_top.sv"
endpackage
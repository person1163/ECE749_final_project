  import uvm_pkg::*;
import decode_in_pkg::*;
import decode_out_pkg::*;
import decode_env_pkg::*;
import decode_test_pkg::*;
  module hvl_top();
  initial begin 
    
     run_test();
  end
  endmodule